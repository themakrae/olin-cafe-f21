module test_edge_detectors